module leading_zero_count(input logic [31:0] src,
                          output logic [4:0] count);
    always_comb begin
        casez(src)
            32'b1???????????????????????????????: count = 5'b00000;
            32'b01??????????????????????????????: count = 5'b00001;
            32'b001?????????????????????????????: count = 5'b00010;
            32'b0001????????????????????????????: count = 5'b00011;
            32'b00001???????????????????????????: count = 5'b00100;
            32'b000001??????????????????????????: count = 5'b00101;
            32'b0000001?????????????????????????: count = 5'b00110;
            32'b00000001????????????????????????: count = 5'b00111;
            32'b000000001???????????????????????: count = 5'b01000;
            32'b0000000001??????????????????????: count = 5'b01001;
            32'b00000000001?????????????????????: count = 5'b01010;
            32'b000000000001????????????????????: count = 5'b01011;
            32'b0000000000001???????????????????: count = 5'b01100;
            32'b00000000000001??????????????????: count = 5'b01101;
            32'b000000000000001?????????????????: count = 5'b01110;
            32'b0000000000000001????????????????: count = 5'b01111;
            32'b00000000000000001???????????????: count = 5'b10000;
            32'b000000000000000001??????????????: count = 5'b10001;
            32'b0000000000000000001?????????????: count = 5'b10010;
            32'b00000000000000000001????????????: count = 5'b10011;
            32'b000000000000000000001???????????: count = 5'b10100;
            32'b0000000000000000000001??????????: count = 5'b10101;
            32'b00000000000000000000001?????????: count = 5'b10110;
            32'b000000000000000000000001????????: count = 5'b10111;
            32'b0000000000000000000000001???????: count = 5'b11000;
            32'b00000000000000000000000001??????: count = 5'b11001;
            32'b000000000000000000000000001?????: count = 5'b11010;
            32'b0000000000000000000000000001????: count = 5'b11011;
            32'b00000000000000000000000000001???: count = 5'b11100;
            32'b000000000000000000000000000001??: count = 5'b11101;
            32'b0000000000000000000000000000001?: count = 5'b11110;
            32'b0000_0000_0000_0000_0000_0000_0000_0001: count = 5'b11111;
        endcase
    end
endmodule